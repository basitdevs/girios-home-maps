<svg width="10" height="2" viewBox="0 0 10 2" fill="none" xmlns="http://www.w3.org/2000/svg">
<line x1="0.186523" y1="0.534607" x2="9.46173" y2="0.534608" stroke="#FAFAFA"/>
</svg>
